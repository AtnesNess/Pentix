120
..........
..........
..........
..........
..........
..........
..........
..........
..........
..........
..........
..........
..........
..........
..........
.....444..
.0.1.4441.
.003345113
.003345107
.003325500